.SUBCKT F0 1 25
* COMMAND  : rffilter.py --g chebyshev_0.2 --n 8 --crystal-mesh --l 69.7e-3 --f 4913.57e3 --bw 2400 --ch 3.66e-12
* TYPE     : chebyshev_0.2
* FILTER   : crystal mesh
* ORDER    : 8
* FREQ     : 4.915464 MHz
* RS       : 1153.1
* RL       : 1153.0
* CH       : 3.6600e-12
* BW       : 2.4000e+03
* QL       : 2048.1
* QU       : inf
* qo       : inf

* ij        q,k           TD0           TDn           CBW           Q,K
* 01     1.3804  366.1625e-06             -    1.7386e+03    2.8272e+03
* 12     0.7225  368.0723e-06    1.4056e-03    1.7341e+03  352.7866e-06
* 23     0.5602  975.2750e-06    2.1627e-03    1.3445e+03  273.5270e-06
* 34     0.5349  771.7423e-06    1.1676e-03    1.2839e+03  261.1882e-06
* 45     0.5298    1.5964e-03    1.5964e-03    1.2714e+03  258.6605e-06
* 56     0.5349    1.1676e-03  771.7246e-06    1.2839e+03  261.1871e-06
* 67     0.5602    2.1627e-03  975.2995e-06    1.3445e+03  273.5273e-06
* 78     0.7225    1.4056e-03  368.0618e-06    1.7341e+03  352.7876e-06
* 89     1.3804             -  366.1709e-06    1.7386e+03    2.8273e+03

* Xtal       Xtal freq     Mesh freq   Mesh offset
* 1          4913570.0     4914792.1        -672.3
* 2          4913570.0     4915464.4          -0.0
* 3          4913570.0     4915239.2        -225.1
* 4          4913570.0     4915202.7        -261.7
* 5          4913570.0     4915202.7        -261.7
* 6          4913570.0     4915239.2        -225.1
* 7          4913570.0     4915464.4          -0.0
* 8          4913570.0     4914792.1        -672.3

* Xtal              LM          LEFF     %LM Shift
* 1        69.7000e-03  105.5531e-03        51.439
* 2        69.7000e-03  105.5531e-03        51.439
* 3        69.7000e-03  105.5531e-03        51.439
* 4        69.7000e-03  105.5531e-03        51.439
* 5        69.7000e-03  105.5531e-03        51.439
* 6        69.7000e-03  105.5531e-03        51.439
* 7        69.7000e-03  105.5531e-03        51.439
* 8        69.7000e-03  105.5531e-03        51.439

* ij              CKij           CTi
* 12       28.1532e-12   36.3110e-12
* 23       36.3111e-12    7.4808e-06
* 34       38.0265e-12  108.4292e-12
* 45       38.3981e-12   93.2885e-12
* 56       38.0267e-12   93.2876e-12
* 67       36.3111e-12  108.4282e-12
* 78       28.1531e-12    1.0697e-03
* 89                 -   36.3111e-12

C1  1    2      15.0527e-15
L2  2    3      69.7000e-03
C3  1    3       3.6600e-12
C4  3    4      36.3110e-12

C5  4    0      28.1532e-12
C6  4    5      15.0527e-15
L7  5    6      69.7000e-03
C8  4    6       3.6600e-12
C9  6    7       7.4808e-06

C10 7    0      36.3111e-12
C11 7    8      15.0527e-15
L12 8    9      69.7000e-03
C13 7    9       3.6600e-12
C14 9    10    108.4292e-12

C15 10   0      38.0265e-12
C16 10   11     15.0527e-15
L17 11   12     69.7000e-03
C18 10   12      3.6600e-12
C19 12   13     93.2885e-12

C20 13   0      38.3981e-12
C21 13   14     15.0527e-15
L22 14   15     69.7000e-03
C23 13   15      3.6600e-12
C24 15   16     93.2876e-12

C25 16   0      38.0267e-12
C26 16   17     15.0527e-15
L27 17   18     69.7000e-03
C28 16   18      3.6600e-12
C29 18   19    108.4282e-12

C30 19   0      36.3111e-12
C31 19   20     15.0527e-15
L32 20   21     69.7000e-03
C33 19   21      3.6600e-12
C34 21   22      1.0697e-03

C35 22   0      28.1531e-12
C36 22   23     15.0527e-15
L37 23   24     69.7000e-03
C38 22   24      3.6600e-12
C39 24   25     36.3111e-12
.ends
.end

