.SUBCKT F1 1 37
* COMMAND  : rffilter.py -g chebyshev_0.1 -bw 2500 -n 12 -l .0155 -crystal -cp 5e-12 -f 8000017.0,7999933.0,7999940.0,7999945.0,7999985.0,7999996.0,8000000.0,7999991.0,7999966.0,7999945.0,7999939.0,8000026.0
* TYPE     : CHEBYSHEV_0.1
* FILTER   : CRYSTAL_MESH
* ORDER    : 12
* FREQ     : 8.001741 MHz
* RS       : 241.8
* RL       : 239.7
* CP       : 5.0000e-12
* BW       : 2.5000e+03
* QL       : 3200.7
* QU       : inf
* qo       : inf

* ij        q,k           TD0           TDn           CBW           Q,K
* 01     1.2010  305.8321e-06             -    2.0816e+03    3.8440e+03
* 12     0.7560  371.0220e-06    2.2617e-03    1.8899e+03  236.1861e-06
* 23     0.5646  854.0891e-06    3.0755e-03    1.4115e+03  176.4021e-06
* 34     0.5322  788.6446e-06    2.0360e-03    1.3304e+03  166.2691e-06
* 45     0.5214    1.4253e-03    2.5726e-03    1.3035e+03  162.8992e-06
* 56     0.5172    1.2131e-03    1.6315e-03    1.2929e+03  161.5746e-06
* 67     0.5160    1.9990e-03    2.0066e-03    1.2900e+03  161.2156e-06
* 78     0.5171    1.6359e-03    1.2101e-03    1.2927e+03  161.5552e-06
* 89     0.5213    2.5635e-03    1.4312e-03    1.3032e+03  162.8616e-06
* 910    0.5320    2.0418e-03  786.8382e-06    1.3299e+03  166.1990e-06
* 1011   0.5642    3.0655e-03  858.3063e-06    1.4104e+03  176.2658e-06
* 1112   0.7538    2.2691e-03  370.3100e-06    1.8846e+03  235.5240e-06
* 1213   1.2101             -  308.1454e-06    2.0660e+03    3.8731e+03

* Xtal    Xtal freq     Mesh freq   Mesh offset   Xtal offset      LM Shift
* 1       8000017.0     8001111.5        -629.2          84.0      19.259 %
* 2       7999933.0     8001739.0          -1.7           0.0      20.337 %
* 3       7999940.0     8001469.7        -271.0           7.0      20.247 %
* 4       7999945.0     8001418.5        -322.2          12.0      20.182 %
* 5       7999985.0     8001435.0        -305.7          52.0      19.668 %
* 6       7999996.0     8001436.6        -304.1          63.0      19.527 %
* 7       8000000.0     8001440.0        -300.7          67.0      19.476 %
* 8       7999991.0     8001439.2        -301.4          58.0      19.591 %
* 9       7999966.0     8001436.4        -304.2          33.0      19.912 %
* 10      7999945.0     8001472.3        -268.3          12.0      20.182 %
* 11      7999939.0     8001740.7          -0.0           6.0      20.259 %
* 12      8000026.0     8001116.5        -624.2          93.0      19.145 %

* ij              CKij            CSi
* 12       90.2069e-12   136.0937e-12
* 23      120.2819e-12    51.2891e-09
* 34      127.6944e-12   313.3347e-12
* 45      130.6506e-12   263.6841e-12
* 56      132.0819e-12   279.1111e-12
* 67      132.4822e-12   280.9150e-12
* 78      132.1684e-12   284.2570e-12
* 89      130.8699e-12   283.2620e-12
* 910     127.9264e-12   279.9100e-12
* 1011    120.4459e-12   316.6422e-12
* 1112     90.5331e-12    12.2375e-06
* 1213               -   137.3105e-12

C1  1    2      25.5345e-15
L2  2    3      15.5000e-03
C3  1    3       5.0000e-12
C4  3    4     136.0937e-12

C5  4    0      90.2069e-12
C6  4    5      25.5350e-15
L7  5    6      15.5000e-03
C8  4    6       5.0000e-12
C9  6    7      51.2891e-09

C10 7    0     120.2819e-12
C11 7    8      25.5350e-15
L12 8    9      15.5000e-03
C13 7    9       5.0000e-12
C14 9    10    313.3347e-12

C15 10   0     127.6944e-12
C16 10   11     25.5349e-15
L17 11   12     15.5000e-03
C18 10   12      5.0000e-12
C19 12   13    263.6841e-12

C20 13   0     130.6506e-12
C21 13   14     25.5347e-15
L22 14   15     15.5000e-03
C23 13   15      5.0000e-12
C24 15   16    279.1111e-12

C25 16   0     132.0819e-12
C26 16   17     25.5346e-15
L27 17   18     15.5000e-03
C28 16   18      5.0000e-12
C29 18   19    280.9150e-12

C30 19   0     132.4822e-12
C31 19   20     25.5346e-15
L32 20   21     15.5000e-03
C33 19   21      5.0000e-12
C34 21   22    284.2570e-12

C35 22   0     132.1684e-12
C36 22   23     25.5346e-15
L37 23   24     15.5000e-03
C38 22   24      5.0000e-12
C39 24   25    283.2620e-12

C40 25   0     130.8699e-12
C41 25   26     25.5348e-15
L42 26   27     15.5000e-03
C43 25   27      5.0000e-12
C44 27   28    279.9100e-12

C45 28   0     127.9264e-12
C46 28   29     25.5349e-15
L47 29   30     15.5000e-03
C48 28   30      5.0000e-12
C49 30   31    316.6422e-12

C50 31   0     120.4459e-12
C51 31   32     25.5350e-15
L52 32   33     15.5000e-03
C53 31   33      5.0000e-12
C54 33   34     12.2375e-06

C55 34   0      90.5331e-12
C56 34   35     25.5344e-15
L57 35   36     15.5000e-03
C58 34   36      5.0000e-12
C59 36   37    137.3105e-12
.ends
.end

