.SUBCKT F1 1 25
* TYPE:   CHEBYSHEV_02
* FILTER: CRYSTAL_MESH
* ORDER:  8
* FREQ:   4.915110 MHz 
* RS:     1060.0
* RL:     1059.7
* BW:     2.4000e+03
* QL:     2047.3
*
* ij    qi,kij           TD0           TDn           CBW
* 01    1.3800  366.0564e-06             -    1.7391e+03
* 12    0.7225  368.1784e-06    1.4056e-03    1.7341e+03
* 23    0.5602  975.0893e-06    2.1630e-03    1.3444e+03
* 34    0.5349  771.9015e-06    1.1676e-03    1.2839e+03
* 45    0.5298    1.5961e-03    1.5965e-03    1.2715e+03
* 56    0.5349    1.1679e-03  771.7423e-06    1.2838e+03
* 67    0.5601    2.1624e-03  975.4158e-06    1.3443e+03
* 78    0.7225    1.4059e-03  368.1121e-06    1.7341e+03
* 89    1.3803             -  366.1380e-06    1.7387e+03
*
C1  1  2    15.0527e-15
L2  2  3    69.7000e-03
C3  1  3     3.6600e-12
C4  3  4    39.5139e-12

C5  4  0    30.6372e-12
C6  4  5    15.0527e-15
L7  5  6    69.7000e-03
C8  4  6     3.6600e-12
C9  6  7   373.8789e-09

C10 7  0    39.5181e-12
C11 7  8    15.0527e-15
L12 8  9    69.7000e-03
C13 7  9     3.6600e-12
C14 9  10  117.9602e-12

C15 10 0    41.3817e-12
C16 10 11   15.0527e-15
L17 11 12   69.7000e-03
C18 10 12    3.6600e-12
C19 12 13  101.5184e-12

C20 13 0    41.7853e-12
C21 13 14   15.0527e-15
L22 14 15   69.7000e-03
C23 13 15    3.6600e-12
C24 15 16  101.4970e-12

C25 16 0    41.3853e-12
C26 16 17   15.0527e-15
L27 17 18   69.7000e-03
C28 16 18    3.6600e-12
C29 18 19  117.8923e-12

C30 19 0    39.5225e-12
C31 19 20   15.0527e-15
L32 20 21   69.7000e-03
C33 19 21    3.6600e-12
C34 21 22  161.8184e-09

C35 22 0    30.6379e-12
C36 22 23   15.0527e-15
L37 23 24   69.7000e-03
C38 22 24    3.6600e-12
C39 24 25   39.5128e-12
.ends
.end
