.SUBCKT F1 1 4 5 8 9 12 13 16 17 20 21 24 25 28 29 32
* COMMAND  : rffilter.py -g chebyshev_0.2 -n 8 -crystal -l 69.7e-3 -f 4913.57e3 -bw 2400 -cp 3.66e-12
* TYPE     : CHEBYSHEV_0.2
* FILTER   : CRYSTAL_MESH
* ORDER    : 8
* FREQ     : 4.915464 MHz
* RS       : 1153.4
* RL       : 1153.2
* BW       : 2.4000e+03
* QL       : 2048.1

* ij    qi,kij           TD0           TDn           CBW
* 01    1.3800  366.0564e-06             -    1.7391e+03
* 12    0.7225  368.1784e-06    1.4056e-03    1.7341e+03
* 23    0.5602  975.0893e-06    2.1630e-03    1.3444e+03
* 34    0.5349  771.9015e-06    1.1676e-03    1.2839e+03
* 45    0.5298    1.5961e-03    1.5965e-03    1.2715e+03
* 56    0.5349    1.1679e-03  771.7423e-06    1.2838e+03
* 67    0.5601    2.1624e-03  975.4158e-06    1.3443e+03
* 78    0.7225    1.4059e-03  368.1121e-06    1.7341e+03
* 89    1.3803             -  366.1380e-06    1.7387e+03

C1  1    2      15.0527e-15
L2  2    3      69.7000e-03
C3  1    3       3.6600e-12
C4  3    4      36.3085e-12

C5  4    0      28.1524e-12
C6  5    6      15.0527e-15
L7  6    7      69.7000e-03
C8  5    7       3.6600e-12
C9  7    8     298.8735e-09

C10 8    0      36.3129e-12
C11 9    10     15.0527e-15
L12 10   11     69.7000e-03
C13 9    11      3.6600e-12
C14 11   12    108.3878e-12

C15 12   0      38.0254e-12
C16 13   14     15.0527e-15
L17 14   15     69.7000e-03
C18 13   15      3.6600e-12
C19 15   16     93.2808e-12

C20 16   0      38.3962e-12
C21 17   18     15.0527e-15
L22 18   19     69.7000e-03
C23 17   19      3.6600e-12
C24 19   20     93.2612e-12

C25 20   0      38.0287e-12
C26 21   22     15.0527e-15
L27 22   23     69.7000e-03
C28 21   23      3.6600e-12
C29 23   24    108.3253e-12

C30 24   0      36.3170e-12
C31 25   26     15.0527e-15
L32 26   27     69.7000e-03
C33 25   27      3.6600e-12
C34 27   28    139.6574e-09

C35 28   0      28.1530e-12
C36 29   30     15.0527e-15
L37 30   31     69.7000e-03
C38 29   31      3.6600e-12
C39 31   32     36.3075e-12
.ends
.end

