.SUBCKT F1 1 25
* COMMAND  : rffilter.py -k chebyshev_0.5 -bw 2500 -n 8 -l 70e-3 -crystal -f 5000.680e3,5000.123e3,4999.670e3,5000.235e3,5000.320e3,4999.895e3,5000.010e3,5000.485e3
* TYPE     : CHEBYSHEV_0.5
* FILTER   : CRYSTAL_MESH
* ORDER    : 8
* FREQ     : 5.001612 MHz
* RS       : 615.9
* RL       : 615.9
* BW       : 2.5000e+03
* QL       : 2000.6
* QU       : inf

* ij       q,k           TD0           TDn           CBW           Q,K
* 01    1.7850  454.5465e-06             -    1.4006e+03    3.5712e+03
* 12    0.6580  329.4960e-06    1.2890e-03    1.6450e+03  328.8940e-06
* 23    0.5330    1.1473e-03    2.4582e-03    1.3325e+03  266.4141e-06
* 34    0.5150  682.4272e-06    1.0554e-03    1.2875e+03  257.4170e-06
* 45    0.5110    1.8509e-03    1.8172e-03    1.2775e+03  255.4177e-06
* 56    0.5150    1.0299e-03  699.3288e-06    1.2875e+03  257.4170e-06
* 67    0.5330    2.5078e-03    1.1306e-03    1.3325e+03  266.4141e-06
* 78    0.6500    1.2635e-03  337.6566e-06    1.6250e+03  324.8953e-06
* 89    1.7850             -  454.5465e-06    1.4006e+03    3.5712e+03

C1  1    2      14.4705e-15
L2  2    3      70.0000e-03
C3  3    4     331.3895e-12

C4  4    0      43.9918e-12
C5  4    5      14.4737e-15
L6  5    6      70.0000e-03
C7  6    7       9.8994e-06

C8  7    0      54.3143e-12
C9  7    8      14.4764e-15
L10 8    9      70.0000e-03
C11 9    10     57.2732e-12

C12 10   0      56.2120e-12
C13 10   11     14.4731e-15
L14 11   12     70.0000e-03
C15 12   13    383.8459e-12

C16 13   0      56.6483e-12
C17 13   14     14.4726e-15
L18 14   15     70.0000e-03
C19 15   16      3.9129e-09

C20 16   0      56.2103e-12
C21 16   17     14.4751e-15
L22 17   18     70.0000e-03
C23 18   19     88.9534e-12

C24 19   0      54.3137e-12
C25 19   20     14.4744e-15
L26 20   21     70.0000e-03
C27 21   22    294.1400e-12

C28 22   0      44.5346e-12
C29 22   23     14.4716e-15
L30 23   24     70.0000e-03
C31 24   25    115.1531e-12
.ends
.end

