.SUBCKT F1 1 5 6 10 11 15 16 20 21 25 26 30 31 35 36 40
* COMMAND  : rffilter.py -g chebyshev_0.2 -n 8 -crystal -l 69.7e-3 -f 4913.57e3 -bw 2400 -cp 3.66e-12 -qu 150000
* TYPE     : CHEBYSHEV_0.2
* FILTER   : CRYSTAL_MESH
* ORDER    : 8
* FREQ     : 4.915464 MHz
* RS       : 1153.4
* RL       : 1153.2
* BW       : 2.4000e+03
* QL       : 2048.1
* QU       : 150000.0

* ij    qi,kij           TD0           TDn           CBW
* 01    1.3800  366.0564e-06             -    1.7391e+03
* 12    0.7225  368.1784e-06    1.4056e-03    1.7341e+03
* 23    0.5602  975.0893e-06    2.1630e-03    1.3444e+03
* 34    0.5349  771.9015e-06    1.1676e-03    1.2839e+03
* 45    0.5298    1.5961e-03    1.5965e-03    1.2715e+03
* 56    0.5349    1.1679e-03  771.7423e-06    1.2838e+03
* 67    0.5601    2.1624e-03  975.4158e-06    1.3443e+03
* 78    0.7225    1.4059e-03  368.1121e-06    1.7341e+03
* 89    1.3803             -  366.1380e-06    1.7387e+03

C1  1    2      15.0527e-15
L2  2    3      69.7000e-03
R3  3    4      14.3511e+00
C4  1    4       3.6600e-12
C5  4    5      36.3097e-12

C6  5    0      28.1527e-12
C7  6    7      15.0527e-15
L8  7    8      69.7000e-03
R9  8    9      14.3511e+00
C10 6    9       3.6600e-12
C11 9    10    362.1959e-09

C12 10   0      36.3134e-12
C13 11   12     15.0527e-15
L14 12   13     69.7000e-03
R15 13   14     14.3511e+00
C16 11   14      3.6600e-12
C17 14   15    108.3959e-12

C18 15   0      38.0259e-12
C19 16   17     15.0527e-15
L20 17   18     69.7000e-03
R21 18   19     14.3511e+00
C22 16   19      3.6600e-12
C23 19   20     93.2870e-12

C24 20   0      38.3967e-12
C25 21   22     15.0527e-15
L26 22   23     69.7000e-03
R27 23   24     14.3511e+00
C28 21   24      3.6600e-12
C29 24   25     93.2674e-12

C30 25   0      38.0291e-12
C31 26   27     15.0527e-15
L32 27   28     69.7000e-03
R33 28   29     14.3511e+00
C34 26   29      3.6600e-12
C35 29   30    108.3335e-12

C36 30   0      36.3174e-12
C37 31   32     15.0527e-15
L38 32   33     69.7000e-03
R39 33   34     14.3511e+00
C40 31   34      3.6600e-12
C41 34   35    152.0826e-09

C42 35   0      28.1533e-12
C43 36   37     15.0527e-15
L44 37   38     69.7000e-03
R45 38   39     14.3511e+00
C46 36   39      3.6600e-12
C47 39   40     36.3087e-12
.ends
.end

