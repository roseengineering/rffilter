.SUBCKT F1 1 49
* COMMAND  : rffilter.py -g chebyshev_0.1 -bw 2500 -n 12 -l .0155 -crystal -cp 5e-12 -qu 120000 -f 8000017.0,7999933.0,7999940.0,7999945.0,7999985.0,7999996.0,8000000.0,7999991.0,7999966.0,7999945.0,7999939.0,8000026.0
* TYPE     : CHEBYSHEV_0.1
* FILTER   : CRYSTAL_MESH
* ORDER    : 12
* FREQ     : 8.001741 MHz
* RS       : 241.8
* RL       : 239.7
* CP       : 5.0000e-12
* BW       : 2.5000e+03
* QL       : 3200.7
* QU       : 120000.0

* ij        q,k           TD0           TDn           CBW           Q,K
* 01     1.2010  305.8321e-06             -    2.0816e+03    3.8440e+03
* 12     0.7560  371.0220e-06    2.2617e-03    1.8899e+03  236.1861e-06
* 23     0.5646  854.0891e-06    3.0755e-03    1.4115e+03  176.4021e-06
* 34     0.5322  788.6446e-06    2.0360e-03    1.3304e+03  166.2691e-06
* 45     0.5214    1.4253e-03    2.5726e-03    1.3035e+03  162.8992e-06
* 56     0.5172    1.2131e-03    1.6315e-03    1.2929e+03  161.5746e-06
* 67     0.5160    1.9990e-03    2.0066e-03    1.2900e+03  161.2156e-06
* 78     0.5171    1.6359e-03    1.2101e-03    1.2927e+03  161.5552e-06
* 89     0.5213    2.5635e-03    1.4312e-03    1.3032e+03  162.8616e-06
* 910    0.5320    2.0418e-03  786.8382e-06    1.3299e+03  166.1990e-06
* 1011   0.5642    3.0655e-03  858.3063e-06    1.4104e+03  176.2658e-06
* 1112   0.7538    2.2691e-03  370.3100e-06    1.8846e+03  235.5240e-06
* 1213   1.2101             -  308.1454e-06    2.0660e+03    3.8731e+03

* Xtal    Xtal freq     Mesh freq   Mesh offset   Xtal offset      LM Shift
* 1       8000017.0     8001111.6        -629.2          84.0       19.259%
* 2       7999933.0     8001739.1          -1.7           0.0       20.336%
* 3       7999940.0     8001469.7        -271.0           7.0       20.246%
* 4       7999945.0     8001418.5        -322.2          12.0       20.182%
* 5       7999985.0     8001435.0        -305.7          52.0       19.668%
* 6       7999996.0     8001436.6        -304.1          63.0       19.527%
* 7       8000000.0     8001440.1        -300.7          67.0       19.476%
* 8       7999991.0     8001439.3        -301.5          58.0       19.591%
* 9       7999966.0     8001436.5        -304.2          33.0       19.911%
* 10      7999945.0     8001472.4        -268.3          12.0       20.182%
* 11      7999939.0     8001740.7          -0.0           6.0       20.259%
* 12      8000026.0     8001116.5        -624.2          93.0       19.145%

* ij              CKij            CSi
* 12       90.2072e-12   136.0932e-12
* 23      120.2823e-12    51.1527e-09
* 34      127.6948e-12   313.3307e-12
* 45      130.6510e-12   263.6813e-12
* 56      132.0823e-12   279.1079e-12
* 67      132.4827e-12   280.9119e-12
* 78      132.1689e-12   284.2538e-12
* 89      130.8704e-12   283.2588e-12
* 910     127.9268e-12   279.9069e-12
* 1011    120.4463e-12   316.6380e-12
* 1112     90.5334e-12     7.4798e-06
* 1213               -   137.3100e-12

C1  1    2      25.5345e-15
L2  2    3      15.5000e-03
R3  3    4       6.4940e+00
C4  1    4       5.0000e-12
C5  4    5     136.0932e-12

C6  5    0      90.2072e-12
C7  5    6      25.5350e-15
L8  6    7      15.5000e-03
R9  7    8       6.4940e+00
C10 5    8       5.0000e-12
C11 8    9      51.1527e-09

C12 9    0     120.2823e-12
C13 9    10     25.5350e-15
L14 10   11     15.5000e-03
R15 11   12      6.4940e+00
C16 9    12      5.0000e-12
C17 12   13    313.3307e-12

C18 13   0     127.6948e-12
C19 13   14     25.5349e-15
L20 14   15     15.5000e-03
R21 15   16      6.4940e+00
C22 13   16      5.0000e-12
C23 16   17    263.6813e-12

C24 17   0     130.6510e-12
C25 17   18     25.5347e-15
L26 18   19     15.5000e-03
R27 19   20      6.4940e+00
C28 17   20      5.0000e-12
C29 20   21    279.1079e-12

C30 21   0     132.0823e-12
C31 21   22     25.5346e-15
L32 22   23     15.5000e-03
R33 23   24      6.4940e+00
C34 21   24      5.0000e-12
C35 24   25    280.9119e-12

C36 25   0     132.4827e-12
C37 25   26     25.5346e-15
L38 26   27     15.5000e-03
R39 27   28      6.4940e+00
C40 25   28      5.0000e-12
C41 28   29    284.2538e-12

C42 29   0     132.1689e-12
C43 29   30     25.5346e-15
L44 30   31     15.5000e-03
R45 31   32      6.4940e+00
C46 29   32      5.0000e-12
C47 32   33    283.2588e-12

C48 33   0     130.8704e-12
C49 33   34     25.5348e-15
L50 34   35     15.5000e-03
R51 35   36      6.4940e+00
C52 33   36      5.0000e-12
C53 36   37    279.9069e-12

C54 37   0     127.9268e-12
C55 37   38     25.5349e-15
L56 38   39     15.5000e-03
R57 39   40      6.4940e+00
C58 37   40      5.0000e-12
C59 40   41    316.6380e-12

C60 41   0     120.4463e-12
C61 41   42     25.5350e-15
L62 42   43     15.5000e-03
R63 43   44      6.4940e+00
C64 41   44      5.0000e-12
C65 44   45      7.4798e-06

C66 45   0      90.5334e-12
C67 45   46     25.5344e-15
L68 46   47     15.5000e-03
R69 47   48      6.4940e+00
C70 45   48      5.0000e-12
C71 48   49    137.3100e-12
.ends
.end

