.SUBCKT F1 1 37
* COMMAND  : rffilter.py -g chebyshev_0.1 -bw 2500 -n 12 -l .0155 -crystal -cp 5e-12 -f 8000017.0,7999966.0,7999940.0,7999945.0,7999985.0,8000000.0,7999996.0,7999991.0,7999939.0,7999933.0,7999945.0,8000026.0
* TYPE     : CHEBYSHEV_0.1
* FILTER   : CRYSTAL_MESH
* ORDER    : 12
* FREQ     : 8.001775 MHz
* RS       : 242.7
* RL       : 240.6
* CP       : 5.0000e-12
* BW       : 2.5000e+03
* QL       : 3200.7
* QU       : inf

* ij        q,k           TD0           TDn           CBW           Q,K
* 01     1.2010  305.8321e-06             -    2.0816e+03    3.8441e+03
* 12     0.7560  371.0220e-06    2.2617e-03    1.8899e+03  236.1850e-06
* 23     0.5646  854.0891e-06    3.0755e-03    1.4115e+03  176.4013e-06
* 34     0.5322  788.6446e-06    2.0360e-03    1.3304e+03  166.2684e-06
* 45     0.5214    1.4253e-03    2.5726e-03    1.3035e+03  162.8985e-06
* 56     0.5172    1.2131e-03    1.6315e-03    1.2929e+03  161.5739e-06
* 67     0.5160    1.9990e-03    2.0066e-03    1.2900e+03  161.2149e-06
* 78     0.5171    1.6359e-03    1.2101e-03    1.2927e+03  161.5545e-06
* 89     0.5213    2.5635e-03    1.4312e-03    1.3032e+03  162.8609e-06
* 910    0.5320    2.0418e-03  786.8382e-06    1.3299e+03  166.1983e-06
* 1011   0.5642    3.0655e-03  858.3063e-06    1.4104e+03  176.2650e-06
* 1112   0.7538    2.2691e-03  370.3100e-06    1.8846e+03  235.5230e-06
* 1213   1.2101             -  308.1454e-06    2.0660e+03    3.8731e+03

* Xtal    Xtal freq     Mesh freq   Mesh offset   Xtal offset      LM Shift
* 1       8000017.0     8001115.7        -659.5          84.0       19.701%
* 2       7999966.0     8001775.2          -0.0          33.0       20.357%
* 3       7999940.0     8001474.6        -300.7           7.0       20.693%
* 4       7999945.0     8001424.6        -350.7          12.0       20.629%
* 5       7999985.0     8001440.8        -334.4          52.0       20.112%
* 6       8000000.0     8001446.2        -329.0          67.0       19.919%
* 7       7999996.0     8001442.2        -333.0          63.0       19.970%
* 8       7999991.0     8001446.3        -328.9          58.0       20.035%
* 9       7999939.0     8001418.8        -356.4           6.0       20.706%
* 10      7999933.0     8001468.5        -306.7           0.0       20.784%
* 11      7999945.0     8001752.7         -22.5          12.0       20.629%
* 12      8000026.0     8001122.0        -653.2          93.0       19.586%

* ij              CKij            CSi
* 12       90.0326e-12   129.3563e-12
* 23      120.0486e-12    13.1039e-06
* 34      127.2212e-12   281.3962e-12
* 45      130.1670e-12   241.4203e-12
* 56      131.6219e-12   254.2288e-12
* 67      131.9927e-12   258.8368e-12
* 78      131.6518e-12   255.6140e-12
* 89      130.1970e-12   258.6378e-12
* 910     127.1859e-12   237.3806e-12
* 1011    119.9609e-12   275.6183e-12
* 1112     90.2273e-12     3.7629e-09
* 1213               -   130.7340e-12

C1  1    2      25.5345e-15
L2  2    3      15.5000e-03
C3  1    3       5.0000e-12
C4  3    4     129.3563e-12

C5  4    0      90.0326e-12
C6  4    5      25.5348e-15
L7  5    6      15.5000e-03
C8  4    6       5.0000e-12
C9  6    7      13.1039e-06

C10 7    0     120.0486e-12
C11 7    8      25.5350e-15
L12 8    9      15.5000e-03
C13 7    9       5.0000e-12
C14 9    10    281.3962e-12

C15 10   0     127.2212e-12
C16 10   11     25.5349e-15
L17 11   12     15.5000e-03
C18 10   12      5.0000e-12
C19 12   13    241.4203e-12

C20 13   0     130.1670e-12
C21 13   14     25.5347e-15
L22 14   15     15.5000e-03
C23 13   15      5.0000e-12
C24 15   16    254.2288e-12

C25 16   0     131.6219e-12
C26 16   17     25.5346e-15
L27 17   18     15.5000e-03
C28 16   18      5.0000e-12
C29 18   19    258.8368e-12

C30 19   0     131.9927e-12
C31 19   20     25.5346e-15
L32 20   21     15.5000e-03
C33 19   21      5.0000e-12
C34 21   22    255.6140e-12

C35 22   0     131.6518e-12
C36 22   23     25.5346e-15
L37 23   24     15.5000e-03
C38 22   24      5.0000e-12
C39 24   25    258.6378e-12

C40 25   0     130.1970e-12
C41 25   26     25.5350e-15
L42 26   27     15.5000e-03
C43 25   27      5.0000e-12
C44 27   28    237.3806e-12

C45 28   0     127.1859e-12
C46 28   29     25.5350e-15
L47 29   30     15.5000e-03
C48 28   30      5.0000e-12
C49 30   31    275.6183e-12

C50 31   0     119.9609e-12
C51 31   32     25.5349e-15
L52 32   33     15.5000e-03
C53 31   33      5.0000e-12
C54 33   34      3.7629e-09

C55 34   0      90.2273e-12
C56 34   35     25.5344e-15
L57 35   36     15.5000e-03
C58 34   36      5.0000e-12
C59 36   37    130.7340e-12
.ends
.end

