.SUBCKT F0 1 33
* COMMAND  : rffilter.py --g chebyshev_0.2 --n 8 --crystal-mesh --l 69.7e-3 --f 4913.57e3 --bw 2400 --ch 3.66e-12 --qu 150000
* TYPE     : chebyshev_0.2
* FILTER   : crystal mesh
* ORDER    : 8
* FREQ     : 4.915464 MHz
* RE1      : 1153.066
* RE2      : 1153.040
* CH       : 3.6600e-12
* BW       : 2.4000e+03
* QL       : 2048.1
* QU       : 150000.0
* qo       : 73.2
* TD21     : 892.0701e-06

* ij        q,k           TD1           TDN           CBW           Q,K      QU/QE>10
* 1      1.3804  366.1625e-06             -    1.7386e+03    2.8272e+03   53.0558e+00
* 12     0.7225  368.0723e-06    1.4056e-03    1.7341e+03  352.7866e-06   52.9180e+00
* 23     0.5602  975.2750e-06    2.1627e-03    1.3445e+03  273.5270e-06   41.0291e+00
* 34     0.5349  771.7423e-06    1.1676e-03    1.2839e+03  261.1882e-06   39.1782e+00
* 45     0.5298    1.5964e-03    1.5964e-03    1.2714e+03  258.6605e-06   38.7991e+00
* 56     0.5349    1.1676e-03  771.7246e-06    1.2839e+03  261.1871e-06   39.1781e+00
* 67     0.5602    2.1627e-03  975.2995e-06    1.3445e+03  273.5273e-06   41.0291e+00
* 78     0.7225    1.4056e-03  368.0618e-06    1.7341e+03  352.7876e-06   52.9181e+00
* 8      1.3804             -  366.1709e-06    1.7386e+03    2.8273e+03   53.0546e+00

* Group Delay for Lossy Q Resonators
* i         q,k           TDn            QU
* 1      1.3804  366.2926e-06  150.0000e+03
* 2      0.7225  367.8102e-06  150.0000e+03
* 3      0.5602  976.6501e-06  150.0000e+03
* 4      0.5349  770.4380e-06  150.0000e+03
* 5      0.5298    1.6015e-03  150.0000e+03
* 6      0.5349    1.1640e-03  150.0000e+03
* 7      0.5602    2.1746e-03  150.0000e+03
* -- reversed --
* i         q,k           TDn            QU
* 8      1.3804  366.3011e-06  150.0000e+03
* 7      0.7225  367.7996e-06  150.0000e+03
* 6      0.5602  976.6748e-06  150.0000e+03
* 5      0.5349  770.4202e-06  150.0000e+03
* 4      0.5298    1.6015e-03  150.0000e+03
* 3      0.5349    1.1640e-03  150.0000e+03
* 2      0.5602    2.1746e-03  150.0000e+03

* Xtal       Xtal freq     Mesh freq   Mesh offset
* 1          4913570.0     4914792.1        -672.3
* 2          4913570.0     4915464.4          -0.0
* 3          4913570.0     4915239.2        -225.1
* 4          4913570.0     4915202.7        -261.7
* 5          4913570.0     4915202.7        -261.7
* 6          4913570.0     4915239.2        -225.1
* 7          4913570.0     4915464.4          -0.0
* 8          4913570.0     4914792.1        -672.3

* Xtal              LM          LEFF     %LM Shift
* 1        69.7000e-03  105.5524e-03        51.438
* 2        69.7000e-03  105.5524e-03        51.438
* 3        69.7000e-03  105.5524e-03        51.438
* 4        69.7000e-03  105.5524e-03        51.438
* 5        69.7000e-03  105.5524e-03        51.438
* 6        69.7000e-03  105.5524e-03        51.438
* 7        69.7000e-03  105.5524e-03        51.438
* 8        69.7000e-03  105.5524e-03        51.438

* ij              CKij           CTi
* 12       28.1534e-12   36.3112e-12
* 23       36.3114e-12    7.5262e-06
* 34       38.0268e-12  108.4299e-12
* 45       38.3984e-12   93.2892e-12
* 56       38.0269e-12   93.2882e-12
* 67       36.3113e-12  108.4289e-12
* 78       28.1533e-12    7.6701e-03
* 89                 -   36.3113e-12

C1  1    2      15.0527e-15
L2  2    3      69.7000e-03
R3  3    4      14.3511e+00
C4  1    4       3.6600e-12
C5  4    5      36.3112e-12

C6  5    0      28.1534e-12
C7  5    6      15.0527e-15
L8  6    7      69.7000e-03
R9  7    8      14.3511e+00
C10 5    8       3.6600e-12
C11 8    9       7.5262e-06

C12 9    0      36.3114e-12
C13 9    10     15.0527e-15
L14 10   11     69.7000e-03
R15 11   12     14.3511e+00
C16 9    12      3.6600e-12
C17 12   13    108.4299e-12

C18 13   0      38.0268e-12
C19 13   14     15.0527e-15
L20 14   15     69.7000e-03
R21 15   16     14.3511e+00
C22 13   16      3.6600e-12
C23 16   17     93.2892e-12

C24 17   0      38.3984e-12
C25 17   18     15.0527e-15
L26 18   19     69.7000e-03
R27 19   20     14.3511e+00
C28 17   20      3.6600e-12
C29 20   21     93.2882e-12

C30 21   0      38.0269e-12
C31 21   22     15.0527e-15
L32 22   23     69.7000e-03
R33 23   24     14.3511e+00
C34 21   24      3.6600e-12
C35 24   25    108.4289e-12

C36 25   0      36.3113e-12
C37 25   26     15.0527e-15
L38 26   27     69.7000e-03
R39 27   28     14.3511e+00
C40 25   28      3.6600e-12
C41 28   29      7.6701e-03

C42 29   0      28.1533e-12
C43 29   30     15.0527e-15
L44 30   31     69.7000e-03
R45 31   32     14.3511e+00
C46 29   32      3.6600e-12
C47 32   33     36.3113e-12
.ends
.end

