.SUBCKT F1 1 4 5 8 9 12 13 16 17 20 21 24 25 28 29 32
* COMMAND  : rffilter.py -k chebyshev_0.1 -n 8 -crystal -l .170 -f 4e6 -bw 500 -cp 2.05e-12 -expose
* TYPE     : CHEBYSHEV_0.1
* FILTER   : CRYSTAL_MESH
* ORDER    : 8
* FREQ     : 4.000330 MHz
* RS       : 459.7
* RL       : 459.7
* CP       : 2.0500e-12
* BW       : 500.0000e+00
* QL       : 8000.7
* QU       : inf

* ij       q,k           TD0           TDn           CBW           Q,K
* 01    1.2510    1.5928e-03             -  399.6803e+00   10.0088e+03
* 12    0.7280    1.9204e-03    7.3284e-03  364.0000e+00   90.9925e-06
* 23    0.5450    4.4349e-03    9.9522e-03  272.5000e+00   68.1194e-06
* 34    0.5160    4.0627e-03    6.1555e-03  258.0000e+00   64.4947e-06
* 45    0.5100    7.3443e-03    7.3443e-03  255.0000e+00   63.7447e-06
* 56    0.5160    6.1555e-03    4.0627e-03  258.0000e+00   64.4947e-06
* 67    0.5450    9.9522e-03    4.4349e-03  272.5000e+00   68.1194e-06
* 78    0.7280    7.3284e-03    1.9204e-03  364.0000e+00   90.9925e-06
* 89    1.2510             -    1.5928e-03  399.6803e+00   10.0088e+03

* Xtal         Mesh       Offset
*    1    4000194.0       -136.3
*    2    4000330.2         -0.0
*    3    4000277.2        -53.0
*    4    4000268.5        -61.8
*    5    4000268.5        -61.8
*    6    4000277.2        -53.0
*    7    4000330.2         -0.0
*    8    4000194.0       -136.3

C1  1    2       9.3126e-15
L2  2    3     170.0000e-03
C3  1    3       2.0500e-12
C4  3    4     126.9354e-12

C5  4    0      95.0313e-12
C6  5    6       9.3126e-15
L7  6    7     170.0000e-03
C8  5    7       2.0500e-12
C9  7    8       2.9216e-06

C10 8    0     126.9409e-12
C11 9    10      9.3126e-15
L12 10   11    170.0000e-03
C13 9    11      2.0500e-12
C14 11   12    326.2975e-12

C15 12   0     134.0752e-12
C16 13   14      9.3126e-15
L17 14   15    170.0000e-03
C18 13   15      2.0500e-12
C19 15   16    280.0655e-12

C20 16   0     135.6526e-12
C21 17   18      9.3126e-15
L22 18   19    170.0000e-03
C23 17   19      2.0500e-12
C24 19   20    280.0655e-12

C25 20   0     134.0752e-12
C26 21   22      9.3126e-15
L27 22   23    170.0000e-03
C28 21   23      2.0500e-12
C29 23   24    326.2975e-12

C30 24   0     126.9409e-12
C31 25   26      9.3126e-15
L32 26   27    170.0000e-03
C33 25   27      2.0500e-12
C34 27   28      2.9216e-06

C35 28   0      95.0313e-12
C36 29   30      9.3126e-15
L37 30   31    170.0000e-03
C38 29   31      2.0500e-12
C39 31   32    126.9354e-12
.ends
.end

