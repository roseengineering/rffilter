.SUBCKT F1 1 25
* COMMAND  : rffilter.py -k chebyshev_0.5 -bw 2500 -n 8 -l 70e-3 -crystal -cp 3.7e-12 -f 5000.680e3,5000.123e3,4999.670e3,5000.235e3,5000.320e3,4999.895e3,5000.010e3,5000.485e3
* TYPE     : CHEBYSHEV_0.5
* FILTER   : CRYSTAL_MESH
* ORDER    : 8
* FREQ     : 5.001933 MHz
* RS       : 810.2
* RL       : 848.6
* CP       : 3.7000e-12
* BW       : 2.5000e+03
* QL       : 2000.8
* QU       : inf

* ij        q,k           TD0           TDn           CBW           Q,K
* 01     1.7850  454.5465e-06             -    1.4006e+03    3.5714e+03
* 12     0.6580  329.4960e-06    1.2579e-03    1.6450e+03  328.8729e-06
* 23     0.5330    1.1473e-03    2.5078e-03    1.3325e+03  266.3970e-06
* 34     0.5150  682.4272e-06    1.0299e-03    1.2875e+03  257.4005e-06
* 45     0.5110    1.8509e-03    1.8509e-03    1.2775e+03  255.4013e-06
* 56     0.5150    1.0299e-03  682.4272e-06    1.2875e+03  257.4005e-06
* 67     0.5330    2.5078e-03    1.1473e-03    1.3325e+03  266.3970e-06
* 78     0.6580    1.2579e-03  329.4960e-06    1.6450e+03  328.8729e-06
* 89     1.7850             -  454.5465e-06    1.4006e+03    3.5714e+03

* Xtal    Xtal freq     Mesh freq   Mesh offset   Xtal offset
* 1       5000680.0     5001720.4        -212.7        1010.0
* 2       5000123.0     5001933.1          -0.0         453.0
* 3       4999670.0     5001420.7        -512.4           0.0
* 4       5000235.0     5001854.0         -79.1         565.0
* 5       5000320.0     5001910.5         -22.6         650.0
* 6       4999895.0     5001586.4        -346.7         225.0
* 7       5000010.0     5001839.8         -93.3         340.0
* 8       5000485.0     5001571.5        -361.6         815.0

* ij               CKij             CSi
* 12       -31.2521e-12   -129.3251e-12
* 23       -34.0134e-12     -4.1971e-06
* 34       -35.6967e-12    -41.7146e-12
* 45       -39.0856e-12   -312.2147e-12
* 56       -37.1512e-12     -1.1170e-09
* 67       -34.5346e-12    -65.3900e-12
* 78       -30.1050e-12   -250.3087e-12
* 89                  -    -72.6241e-12

C1  1    2      14.4705e-15
L2  2    3      70.0000e-03
C3  1    3       3.7000e-12
C4  3    4     129.3251e-12

C5  4    0      31.2521e-12
C6  4    5      14.4737e-15
L7  5    6      70.0000e-03
C8  4    6       3.7000e-12
C9  6    7       4.1971e-06

C10 7    0      34.0134e-12
C11 7    8      14.4764e-15
L12 8    9      70.0000e-03
C13 7    9       3.7000e-12
C14 9    10     41.7146e-12

C15 10   0      35.6967e-12
C16 10   11     14.4731e-15
L17 11   12     70.0000e-03
C18 10   12      3.7000e-12
C19 12   13    312.2147e-12

C20 13   0      39.0856e-12
C21 13   14     14.4726e-15
L22 14   15     70.0000e-03
C23 13   15      3.7000e-12
C24 15   16      1.1170e-09

C25 16   0      37.1512e-12
C26 16   17     14.4751e-15
L27 17   18     70.0000e-03
C28 16   18      3.7000e-12
C29 18   19     65.3900e-12

C30 19   0      34.5346e-12
C31 19   20     14.4744e-15
L32 20   21     70.0000e-03
C33 19   21      3.7000e-12
C34 21   22    250.3087e-12

C35 22   0      30.1050e-12
C36 22   23     14.4716e-15
L37 23   24     70.0000e-03
C38 22   24      3.7000e-12
C39 24   25     72.6241e-12
.ends
.end

