.SUBCKT F1 1 25
* COMMAND  : rffilter.py -g chebyshev_0.2 -n 8 -crystal -l 69.7e-3 -f 4913.57e3 -bw 2400 -cp 3.66e-12
* TYPE     : CHEBYSHEV_0.2
* FILTER   : CRYSTAL_MESH
* ORDER    : 8
* FREQ     : 4.915464 MHz
* RS       : 1153.4
* RL       : 1153.1
* CP       : 3.6600e-12
* BW       : 2.4000e+03
* QL       : 2048.1
* QU       : inf

* ij       q,k           TD0           TDn           CBW           Q,K
* 01    1.3800  366.0564e-06             -    1.7391e+03    2.8264e+03
* 12    0.7225  368.1784e-06    1.4056e-03    1.7341e+03  352.7869e-06
* 23    0.5602  975.0893e-06    2.1630e-03    1.3444e+03  273.5055e-06
* 34    0.5349  771.9015e-06    1.1676e-03    1.2839e+03  261.1881e-06
* 45    0.5298    1.5961e-03    1.5965e-03    1.2715e+03  258.6656e-06
* 56    0.5349    1.1679e-03  771.7423e-06    1.2838e+03  261.1657e-06
* 67    0.5601    2.1624e-03  975.4158e-06    1.3443e+03  273.4751e-06
* 78    0.7225    1.4059e-03  368.1121e-06    1.7341e+03  352.7793e-06
* 89    1.3803             -  366.1380e-06    1.7387e+03    2.8270e+03

* Xtal         Mesh       Offset
*    1    4914792.0       -672.3
*    2    4915464.3         -0.0
*    3    4915239.1       -225.1
*    4    4915202.7       -261.6
*    5    4915202.6       -261.7
*    6    4915239.0       -225.3
*    7    4915464.2         -0.1
*    8    4914792.0       -672.3

C1  1    2      15.0527e-15
L2  2    3      69.7000e-03
C3  1    3       3.6600e-12
C4  3    4      36.3145e-12

C5  4    0      28.1538e-12
C6  4    5      15.0527e-15
L7  5    6      69.7000e-03
C8  4    6       3.6600e-12
C9  6    7       5.8570e-06

C10 7    0      36.3147e-12
C11 7    8      15.0527e-15
L12 8    9      69.7000e-03
C13 7    9       3.6600e-12
C14 9    10    108.4305e-12

C15 10   0      38.0273e-12
C16 10   11     15.0527e-15
L17 11   12     69.7000e-03
C18 10   12      3.6600e-12
C19 12   13     93.3131e-12

C20 13   0      38.3981e-12
C21 13   14     15.0527e-15
L22 14   15     69.7000e-03
C23 13   15      3.6600e-12
C24 15   16     93.2934e-12

C25 16   0      38.0306e-12
C26 16   17     15.0527e-15
L27 17   18     69.7000e-03
C28 16   18      3.6600e-12
C29 18   19    108.3680e-12

C30 19   0      36.3188e-12
C31 19   20     15.0527e-15
L32 20   21     69.7000e-03
C33 19   21      3.6600e-12
C34 21   22    250.9392e-09

C35 22   0      28.1544e-12
C36 22   23     15.0527e-15
L37 23   24     69.7000e-03
C38 22   24      3.6600e-12
C39 24   25     36.3135e-12
.ends
.end

