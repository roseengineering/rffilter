.SUBCKT F0 1 17
* COMMAND  : rffilter.py -g butterworth -mesh -f 10e6 -bw 400e3 -n 8
* TYPE     : BUTTERWORTH
* FILTER   : MESH
* ORDER    : 8
* FREQ     : 10.000000 MHz
* RS       : 50.0
* RL       : 50.0
* BW       : 400.0000e+03
* QL       : 25.0
* QU       : inf
* qo       : inf

* ij        q,k           TD0           TDn           CBW           Q,K
* 01     0.3902  621.0226e-09             -    1.0251e+06    9.7550e+00
* 12     1.5187    1.7684e-06    8.1580e-06  607.4909e+03   60.7491e-03
* 23     0.7357    3.2676e-06    8.1580e-06  294.2730e+03   29.4273e-03
* 34     0.5537    4.8904e-06    7.5369e-06  221.4735e+03   22.1473e-03
* 45     0.5098    6.3896e-06    6.3896e-06  203.9152e+03   20.3915e-03
* 56     0.5537    7.5369e-06    4.8904e-06  221.4735e+03   22.1473e-03
* 67     0.7357    8.1580e-06    3.2676e-06  294.2730e+03   29.4273e-03
* 78     1.5187    8.1580e-06    1.7684e-06  607.4909e+03   60.7491e-03
* 89     0.3902             -  621.0226e-09    1.0251e+06    9.7550e+00

L1  1    2       7.7628e-06
C2  2    3      34.7409e-12

C3  3    0     537.1345e-12
L4  3    4       7.7628e-06
C5  4    5      35.8646e-12

C6  5    0       1.1088e-09
L7  5    6       7.7628e-06
C8  6    7      34.4049e-12

C9  7    0       1.4733e-09
L10 7    8       7.7628e-06
C11 8    9      34.0802e-12

C12 9    0       1.6002e-09
L13 9    10      7.7628e-06
C14 10   11     34.0802e-12

C15 11   0       1.4733e-09
L16 11   12      7.7628e-06
C17 12   13     34.4049e-12

C18 13   0       1.1088e-09
L19 13   14      7.7628e-06
C20 14   15     35.8646e-12

C21 15   0     537.1345e-12
L22 15   16      7.7628e-06
C23 16   17     34.7409e-12
.ends
.end

