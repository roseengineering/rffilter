.SUBCKT F1 1 33
* COMMAND  : rffilter.py -g chebyshev_0.2 -n 8 -crystal -l 69.7e-3 -f 4913.57e3 -bw 2400 -cp 3.66e-12 -qu 150000
* TYPE     : CHEBYSHEV_0.2
* FILTER   : CRYSTAL_MESH
* ORDER    : 8
* FREQ     : 4.915464 MHz
* RS       : 1153.1
* RL       : 1153.1
* CP       : 3.6600e-12
* BW       : 2.4000e+03
* QL       : 2048.1
* QU       : 150000.0
* qo       : 73.2

* ij        q,k           TD0           TDn           CBW           Q,K
* 01     1.3804  366.1625e-06             -    1.7386e+03    2.8272e+03
* 12     0.7225  368.0723e-06    1.4057e-03    1.7341e+03  352.7866e-06
* 23     0.5602  975.2750e-06    2.1625e-03    1.3445e+03  273.5270e-06
* 34     0.5349  771.7423e-06    1.1677e-03    1.2839e+03  261.1882e-06
* 45     0.5298    1.5964e-03    1.5962e-03    1.2714e+03  258.6605e-06
* 56     0.5349    1.1676e-03  771.7940e-06    1.2839e+03  261.1871e-06
* 67     0.5602    2.1627e-03  975.2117e-06    1.3445e+03  273.5273e-06
* 78     0.7225    1.4056e-03  368.0949e-06    1.7341e+03  352.7876e-06
* 89     1.3803             -  366.1380e-06    1.7387e+03    2.8270e+03

* Xtal    Xtal freq     Mesh freq   Mesh offset   Xtal offset      LM Shift
* 1       4913570.0     4914792.1        -672.3           0.0      51.439 %
* 2       4913570.0     4915464.4          -0.0           0.0      51.439 %
* 3       4913570.0     4915239.3        -225.1           0.0      51.439 %
* 4       4913570.0     4915202.7        -261.7           0.0      51.439 %
* 5       4913570.0     4915202.7        -261.7           0.0      51.439 %
* 6       4913570.0     4915239.3        -225.1           0.0      51.439 %
* 7       4913570.0     4915464.4          -0.0           0.0      51.439 %
* 8       4913570.0     4914792.1        -672.3           0.0      51.439 %

* ij              CKij            CSi
* 12       28.1533e-12    36.3108e-12
* 23       36.3113e-12     2.4856e-06
* 34       38.0267e-12   108.4264e-12
* 45       38.3983e-12    93.2866e-12
* 56       38.0268e-12    93.2856e-12
* 67       36.3112e-12   108.4255e-12
* 78       28.1533e-12     3.7094e-06
* 89                 -    36.3109e-12

C1  1    2      15.0527e-15
L2  2    3      69.7000e-03
R3  3    4      14.3511e+00
C4  1    4       3.6600e-12
C5  4    5      36.3108e-12

C6  5    0      28.1533e-12
C7  5    6      15.0527e-15
L8  6    7      69.7000e-03
R9  7    8      14.3511e+00
C10 5    8       3.6600e-12
C11 8    9       2.4856e-06

C12 9    0      36.3113e-12
C13 9    10     15.0527e-15
L14 10   11     69.7000e-03
R15 11   12     14.3511e+00
C16 9    12      3.6600e-12
C17 12   13    108.4264e-12

C18 13   0      38.0267e-12
C19 13   14     15.0527e-15
L20 14   15     69.7000e-03
R21 15   16     14.3511e+00
C22 13   16      3.6600e-12
C23 16   17     93.2866e-12

C24 17   0      38.3983e-12
C25 17   18     15.0527e-15
L26 18   19     69.7000e-03
R27 19   20     14.3511e+00
C28 17   20      3.6600e-12
C29 20   21     93.2856e-12

C30 21   0      38.0268e-12
C31 21   22     15.0527e-15
L32 22   23     69.7000e-03
R33 23   24     14.3511e+00
C34 21   24      3.6600e-12
C35 24   25    108.4255e-12

C36 25   0      36.3112e-12
C37 25   26     15.0527e-15
L38 26   27     69.7000e-03
R39 27   28     14.3511e+00
C40 25   28      3.6600e-12
C41 28   29      3.7094e-06

C42 29   0      28.1533e-12
C43 29   30     15.0527e-15
L44 30   31     69.7000e-03
R45 31   32     14.3511e+00
C46 29   32      3.6600e-12
C47 32   33     36.3109e-12
.ends
.end

