.SUBCKT F1 1 4
* COMMAND  : rffilter.py -g butterworth -lowpass -f 10e6 -n 5
* TYPE     : BUTTERWORTH
* FILTER   : LOWPASS
* ORDER    : 5
* FREQ     : 10.000000 MHz
* RS       : 50.0
* RL       : 50.0
L1  1    2     491.8126e-09

C2  2    0     515.0349e-12
L3  2    3       1.5915e-06

C4  3    0     515.0349e-12
L5  3    4     491.8126e-09
.ends
.end

.SUBCKT F1 1 3
* COMMAND  : rffilter.py -g butterworth -lowpass -f 10e6 -n 5
* TYPE     : BUTTERWORTH
* FILTER   : LOWPASS
* ORDER    : 5
* FREQ     : 10.000000 MHz
* RS       : 50.0
* RL       : 50.0
C1  1    0     196.7251e-12
L2  1    2       1.2876e-06

C3  2    0     636.6198e-12
L4  2    3       1.2876e-06

C5  3    0     196.7251e-12
.ends
.end

