.SUBCKT F1 1 33
* TYPE:   CHEBYSHEV_02
* FILTER: CRYSTAL_MESH
* ORDER:  8
* FREQ:   4.915110 MHz 
* RS:     1060.0
* RL:     1059.7
* BW:     2.4000e+03
* QL:     2047.3
* QU:     150000.0
*
* ij    qi,kij           TD0           TDn           CBW
* 01    1.3800  366.0564e-06             -    1.7391e+03
* 12    0.7225  368.1784e-06    1.4056e-03    1.7341e+03
* 23    0.5602  975.0893e-06    2.1630e-03    1.3444e+03
* 34    0.5349  771.9015e-06    1.1676e-03    1.2839e+03
* 45    0.5298    1.5961e-03    1.5965e-03    1.2715e+03
* 56    0.5349    1.1679e-03  771.7423e-06    1.2838e+03
* 67    0.5601    2.1624e-03  975.4158e-06    1.3443e+03
* 78    0.7225    1.4059e-03  368.1121e-06    1.7341e+03
* 89    1.3803             -  366.1380e-06    1.7387e+03
*
C1  1  2    15.0527e-15
L2  2  3    69.7000e-03
R3  3  4    14.3456e+00
C4  1  4     3.6600e-12
C5  4  5    39.5144e-12

C6  5  0    30.6376e-12
C7  5  6    15.0527e-15
L8  6  7    69.7000e-03
R9  7  8    14.3456e+00
C10 5  8     3.6600e-12
C11 8  9   373.8830e-09

C12 9  0    39.5185e-12
C13 9  10   15.0527e-15
L14 10 11   69.7000e-03
R15 11 12   14.3456e+00
C16 9  12    3.6600e-12
C17 12 13  117.9615e-12

C18 13 0    41.3822e-12
C19 13 14   15.0527e-15
L20 14 15   69.7000e-03
R21 15 16   14.3456e+00
C22 13 16    3.6600e-12
C23 16 17  101.5196e-12

C24 17 0    41.7858e-12
C25 17 18   15.0527e-15
L26 18 19   69.7000e-03
R27 19 20   14.3456e+00
C28 17 20    3.6600e-12
C29 20 21  101.4981e-12

C30 21 0    41.3858e-12
C31 21 22   15.0527e-15
L32 22 23   69.7000e-03
R33 23 24   14.3456e+00
C34 21 24    3.6600e-12
C35 24 25  117.8936e-12

C36 25 0    39.5229e-12
C37 25 26   15.0527e-15
L38 26 27   69.7000e-03
R39 27 28   14.3456e+00
C40 25 28    3.6600e-12
C41 28 29  161.8202e-09

C42 29 0    30.6382e-12
C43 29 30   15.0527e-15
L44 30 31   69.7000e-03
R45 31 32   14.3456e+00
C46 29 32    3.6600e-12
C47 32 33   39.5133e-12
.ends
.end
