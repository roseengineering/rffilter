.SUBCKT F1 1 2 3 4 5
* COMMAND  : rffilter.py -g butterworth -nodal -f 10e6 -bw 400e3 -n 5 -qu 2000
* TYPE     : BUTTERWORTH
* FILTER   : NODAL
* ORDER    : 5
* FREQ     : 10.000000 MHz
* RS       : 50.0
* RL       : 50.0
* BW       : 400.0000e+03
* QL       : 25.0
* QU       : 2000.0

* ij    qi,kij           TD0           TDn           CBW
* 01    0.6180  983.6253e-09             -  647.2178e+03
* 12    1.0000    2.5752e-06    5.1503e-06  400.0018e+03
* 23    0.5559    4.1667e-06    5.1503e-06  222.3575e+03
* 34    0.5559    5.1503e-06    4.1667e-06  222.3575e+03
* 45    1.0000    5.1503e-06    2.5752e-06  400.0018e+03
* 56    0.6180             -  983.6253e-09  647.2178e+03

L1  1    1001   51.5040e-09
R1  1001 0       1.6180e-03
C2  1    0       4.7214e-09
C3  1    2     196.7259e-12

L4  2    1004   51.5040e-09
R4  1004 0       1.6180e-03
C5  2    0       4.6120e-09
C6  2    3     109.3582e-12

L7  3    1007   51.5040e-09
R7  1007 0       1.6180e-03
C8  3    0       4.6994e-09
C9  3    4     109.3582e-12

L10 4    1010   51.5040e-09
R10 1010 0       1.6180e-03
C11 4    0       4.6120e-09
C12 4    5     196.7259e-12

L13 5    1013   51.5040e-09
R13 1013 0       1.6180e-03
C14 5    0       4.7214e-09
.ends
.end

