.SUBCKT F1 1 4 5 8 9 12 13 16 17 20 21 24 25 28 29 32
* COMMAND  : rffilter.py -g chebyshev_0.01 -n 8 -crystal -l .170 -f 4e6 -bw 500 -expose
* TYPE     : CHEBYSHEV_0.01
* FILTER   : CRYSTAL_MESH
* ORDER    : 8
* FREQ     : 4.000392 MHz
* RS       : 661.5
* RL       : 661.5
* BW       : 500.0000e+00
* QL       : 8000.8

* ij    qi,kij           TD0           TDn           CBW
* 01    0.8073    1.0279e-03             -  619.3484e+00
* 12    0.9363    1.7991e-03    6.9373e-03  468.1461e+00
* 23    0.6302    3.2968e-03    7.6358e-03  315.0976e+00
* 34    0.5774    3.9419e-03    6.0035e-03  288.7182e+00
* 45    0.5663    5.6561e-03    5.6555e-03  283.1328e+00
* 56    0.5773    6.0033e-03    3.9422e-03  288.6748e+00
* 67    0.6302    7.6360e-03    3.2968e-03  315.1239e+00
* 78    0.9364    6.9371e-03    1.7987e-03  468.2032e+00
* 89    0.8073             -    1.0278e-03  619.3755e+00

C1  1    2       9.3126e-15
L2  2    3     170.0000e-03
C3  3    4     118.1680e-12

C4  4    0      79.5701e-12
C5  5    6       9.3126e-15
L6  6    7     170.0000e-03
C7  7    8     275.5257e-09

C8  8    0     118.2187e-12
C9  9    10      9.3126e-15
L10 10   11    170.0000e-03
C11 11   12    207.4503e-12

C12 12   0     129.0201e-12
C13 13   14      9.3126e-15
L14 14   15    170.0000e-03
C15 15   16    176.1017e-12

C16 16   0     131.5652e-12
C17 17   18      9.3126e-15
L18 18   19    170.0000e-03
C19 19   20    176.0656e-12

C20 20   0     129.0394e-12
C21 21   22      9.3126e-15
L22 22   23    170.0000e-03
C23 23   24    207.4306e-12

C24 24   0     118.2088e-12
C25 25   26      9.3126e-15
L26 26   27    170.0000e-03
C27 27   28    718.8797e-09

C28 28   0      79.5604e-12
C29 29   30      9.3126e-15
L30 30   31    170.0000e-03
C31 31   32    118.1894e-12
.ends
.end

