.SUBCKT F0 1 37
* COMMAND  : rffilter.py --g chebyshev_0.1 --bw 2500 --n 12 --l .0155 --crystal-mesh --ch 5e-12 --f 8000017.0,7999933.0,7999940.0,7999945.0,7999985.0,7999996.0,8000000.0,7999991.0,7999966.0,7999945.0,7999939.0,8000026.0
* TYPE     : chebyshev_0.1
* FILTER   : crystal mesh
* ORDER    : 12
* FREQ     : 8.001743 MHz
* RE1      : 240.921
* RE2      : 240.691
* CH       : 5.0000e-12
* BW       : 2.5000e+03
* QL       : 3200.7
* QU       : inf
* qo       : inf
* SUM(g1-n): 20.9529e+00
* TD21     : 1.3339e-03

* ij        q,k           TD1           TDN           CBW           Q,K      QU/QE>10
* 1      1.2055  306.9781e-06             -    2.0738e+03    3.8584e+03             -
* 12     0.7550  370.6146e-06    2.2652e-03    1.8874e+03  235.8743e-06             -
* 23     0.5644  856.1517e-06    3.0704e-03    1.4111e+03  176.3516e-06             -
* 34     0.5321  787.7278e-06    2.0388e-03    1.3301e+03  166.2316e-06             -
* 45     0.5213    1.4281e-03    2.5681e-03    1.3033e+03  162.8824e-06             -
* 56     0.5172    1.2116e-03    1.6336e-03    1.2929e+03  161.5758e-06             -
* 67     0.5160    2.0027e-03    2.0027e-03    1.2900e+03  161.2173e-06             -
* 78     0.5172    1.6336e-03    1.2116e-03    1.2929e+03  161.5769e-06             -
* 89     0.5214    2.5680e-03    1.4282e-03    1.3034e+03  162.8889e-06             -
* 910    0.5321    2.0388e-03  787.6913e-06    1.3302e+03  166.2327e-06             -
* 1011   0.5644    3.0703e-03  856.1785e-06    1.4111e+03  176.3492e-06             -
* 1112   0.7550    2.2653e-03  370.6053e-06    1.8874e+03  235.8779e-06             -
* 12     1.2055             -  306.9762e-06    2.0738e+03    3.8584e+03             -

* Xtal       Xtal freq     Mesh freq   Mesh offset
* 1          8000017.0     8001110.6        -632.2
* 2          7999933.0     8001738.0          -4.8
* 3          7999940.0     8001469.7        -273.1
* 4          7999945.0     8001418.6        -324.2
* 5          7999985.0     8001435.3        -307.5
* 6          7999996.0     8001436.9        -305.9
* 7          8000000.0     8001440.5        -302.3
* 8          7999991.0     8001439.8        -303.0
* 9          7999966.0     8001437.1        -305.7
* 10         7999945.0     8001473.2        -269.6
* 11         7999939.0     8001742.8          -0.0
* 12         8000026.0     8001118.3        -624.5

* Xtal              LM          LEFF     %LM Shift
* 1        15.5000e-03   18.4894e-03        19.286
* 2        15.5000e-03   18.6564e-03        20.364
* 3        15.5000e-03   18.6424e-03        20.274
* 4        15.5000e-03   18.6324e-03        20.209
* 5        15.5000e-03   18.5528e-03        19.695
* 6        15.5000e-03   18.5309e-03        19.554
* 7        15.5000e-03   18.5230e-03        19.503
* 8        15.5000e-03   18.5408e-03        19.618
* 9        15.5000e-03   18.5905e-03        19.939
* 10       15.5000e-03   18.6324e-03        20.209
* 11       15.5000e-03   18.6444e-03        20.287
* 12       15.5000e-03   18.4716e-03        19.172

* ij              CKij           CTi
* 12       90.3056e-12  135.4164e-12
* 23      120.2890e-12   17.5537e-09
* 34      127.6942e-12  310.8688e-12
* 45      130.6345e-12  262.0353e-12
* 56      132.0511e-12  277.4077e-12
* 67      132.4509e-12  279.2575e-12
* 78      132.1208e-12  282.6373e-12
* 89      130.8184e-12  281.7490e-12
* 910     127.8715e-12  278.4762e-12
* 1011    120.3617e-12  315.0808e-12
* 1112     90.3768e-12   35.5013e-03
* 1213               -  137.2069e-12

C1  1    2      25.5345e-15
L2  2    3      15.5000e-03
C3  1    3       5.0000e-12
C4  3    4     135.4164e-12

C5  4    0      90.3056e-12
C6  4    5      25.5350e-15
L7  5    6      15.5000e-03
C8  4    6       5.0000e-12
C9  6    7      17.5537e-09

C10 7    0     120.2890e-12
C11 7    8      25.5350e-15
L12 8    9      15.5000e-03
C13 7    9       5.0000e-12
C14 9    10    310.8688e-12

C15 10   0     127.6942e-12
C16 10   11     25.5349e-15
L17 11   12     15.5000e-03
C18 10   12      5.0000e-12
C19 12   13    262.0353e-12

C20 13   0     130.6345e-12
C21 13   14     25.5347e-15
L22 14   15     15.5000e-03
C23 13   15      5.0000e-12
C24 15   16    277.4077e-12

C25 16   0     132.0511e-12
C26 16   17     25.5346e-15
L27 17   18     15.5000e-03
C28 16   18      5.0000e-12
C29 18   19    279.2575e-12

C30 19   0     132.4509e-12
C31 19   20     25.5346e-15
L32 20   21     15.5000e-03
C33 19   21      5.0000e-12
C34 21   22    282.6373e-12

C35 22   0     132.1208e-12
C36 22   23     25.5346e-15
L37 23   24     15.5000e-03
C38 22   24      5.0000e-12
C39 24   25    281.7490e-12

C40 25   0     130.8184e-12
C41 25   26     25.5348e-15
L42 26   27     15.5000e-03
C43 25   27      5.0000e-12
C44 27   28    278.4762e-12

C45 28   0     127.8715e-12
C46 28   29     25.5349e-15
L47 29   30     15.5000e-03
C48 28   30      5.0000e-12
C49 30   31    315.0808e-12

C50 31   0     120.3617e-12
C51 31   32     25.5350e-15
L52 32   33     15.5000e-03
C53 31   33      5.0000e-12
C54 33   34     35.5013e-03

C55 34   0      90.3768e-12
C56 34   35     25.5344e-15
L57 35   36     15.5000e-03
C58 34   36      5.0000e-12
C59 36   37    137.2069e-12
.ends
.end

