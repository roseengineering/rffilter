.SUBCKT F0 1 37
* COMMAND  : rffilter.py --g chebyshev_0.1 --bw 2500 --n 12 --l .0155 --crystal-mesh --ch 5e-12 --f 8000017.0,7999966.0,7999940.0,7999945.0,7999985.0,8000000.0,7999996.0,7999991.0,7999939.0,7999933.0,7999945.0,8000026.0
* TYPE     : chebyshev_0.1
* FILTER   : crystal mesh
* ORDER    : 12
* FREQ     : 8.001773 MHz
* RE1      : 241.7
* RE2      : 241.5
* CH       : 5.0000e-12
* BW       : 2.5000e+03
* QL       : 3200.7
* QU       : inf
* qo       : inf

* ij        q,k           TD1           TDN           CBW           Q,K      QE/QU<.1
* 1      1.2055  306.9781e-06             -    2.0738e+03    3.8585e+03             -
* 12     0.7550  370.6146e-06    2.2652e-03    1.8874e+03  235.8734e-06             -
* 23     0.5644  856.1517e-06    3.0704e-03    1.4111e+03  176.3509e-06             -
* 34     0.5321  787.7278e-06    2.0388e-03    1.3301e+03  166.2310e-06             -
* 45     0.5213    1.4281e-03    2.5681e-03    1.3033e+03  162.8818e-06             -
* 56     0.5172    1.2116e-03    1.6336e-03    1.2929e+03  161.5752e-06             -
* 67     0.5160    2.0027e-03    2.0027e-03    1.2900e+03  161.2167e-06             -
* 78     0.5172    1.6336e-03    1.2116e-03    1.2929e+03  161.5762e-06             -
* 89     0.5214    2.5680e-03    1.4282e-03    1.3034e+03  162.8883e-06             -
* 910    0.5321    2.0388e-03  787.6913e-06    1.3302e+03  166.2321e-06             -
* 1011   0.5644    3.0703e-03  856.1785e-06    1.4111e+03  176.3485e-06             -
* 1112   0.7550    2.2653e-03  370.6053e-06    1.8874e+03  235.8770e-06             -
* 12     1.2055             -  306.9762e-06    2.0738e+03    3.8584e+03             -

* Xtal       Xtal freq     Mesh freq   Mesh offset
* 1          8000017.0     8001114.2        -659.3
* 2          7999966.0     8001773.5          -0.0
* 3          7999940.0     8001473.9        -299.6
* 4          7999945.0     8001424.0        -349.4
* 5          7999985.0     8001440.4        -333.0
* 6          8000000.0     8001445.9        -327.5
* 7          7999996.0     8001442.0        -331.4
* 8          7999991.0     8001446.2        -327.3
* 9          7999939.0     8001418.8        -354.7
* 10         7999933.0     8001468.6        -304.8
* 11         7999945.0     8001754.2         -19.3
* 12         8000026.0     8001123.2        -650.3

* Xtal              LM          LEFF     %LM Shift
* 1        15.5000e-03   18.5501e-03        19.678
* 2        15.5000e-03   18.6518e-03        20.334
* 3        15.5000e-03   18.7039e-03        20.670
* 4        15.5000e-03   18.6939e-03        20.606
* 5        15.5000e-03   18.6138e-03        20.089
* 6        15.5000e-03   18.5839e-03        19.896
* 7        15.5000e-03   18.5919e-03        19.948
* 8        15.5000e-03   18.6018e-03        20.012
* 9        15.5000e-03   18.7059e-03        20.683
* 10       15.5000e-03   18.7180e-03        20.761
* 11       15.5000e-03   18.6939e-03        20.606
* 12       15.5000e-03   18.5323e-03        19.563

* ij              CKij           CTi
* 12       90.1686e-12  129.4220e-12
* 23      120.1057e-12  295.9772e-03
* 34      127.2740e-12  282.4796e-12
* 45      130.2051e-12  242.3174e-12
* 56      131.6458e-12  255.3407e-12
* 67      132.0163e-12  260.0475e-12
* 78      131.6590e-12  256.8588e-12
* 89      130.1998e-12  259.9932e-12
* 910     127.1843e-12  238.5581e-12
* 1011    119.9269e-12  277.4025e-12
* 1112     90.1090e-12    4.3862e-09
* 1213               -  131.3387e-12

C1  1    2      25.5345e-15
L2  2    3      15.5000e-03
C3  1    3       5.0000e-12
C4  3    4     129.4220e-12

C5  4    0      90.1686e-12
C6  4    5      25.5348e-15
L7  5    6      15.5000e-03
C8  4    6       5.0000e-12
C9  6    7     295.9772e-03

C10 7    0     120.1057e-12
C11 7    8      25.5350e-15
L12 8    9      15.5000e-03
C13 7    9       5.0000e-12
C14 9    10    282.4796e-12

C15 10   0     127.2740e-12
C16 10   11     25.5349e-15
L17 11   12     15.5000e-03
C18 10   12      5.0000e-12
C19 12   13    242.3174e-12

C20 13   0     130.2051e-12
C21 13   14     25.5347e-15
L22 14   15     15.5000e-03
C23 13   15      5.0000e-12
C24 15   16    255.3407e-12

C25 16   0     131.6458e-12
C26 16   17     25.5346e-15
L27 17   18     15.5000e-03
C28 16   18      5.0000e-12
C29 18   19    260.0475e-12

C30 19   0     132.0163e-12
C31 19   20     25.5346e-15
L32 20   21     15.5000e-03
C33 19   21      5.0000e-12
C34 21   22    256.8588e-12

C35 22   0     131.6590e-12
C36 22   23     25.5346e-15
L37 23   24     15.5000e-03
C38 22   24      5.0000e-12
C39 24   25    259.9932e-12

C40 25   0     130.1998e-12
C41 25   26     25.5350e-15
L42 26   27     15.5000e-03
C43 25   27      5.0000e-12
C44 27   28    238.5581e-12

C45 28   0     127.1843e-12
C46 28   29     25.5350e-15
L47 29   30     15.5000e-03
C48 28   30      5.0000e-12
C49 30   31    277.4025e-12

C50 31   0     119.9269e-12
C51 31   32     25.5349e-15
L52 32   33     15.5000e-03
C53 31   33      5.0000e-12
C54 33   34      4.3862e-09

C55 34   0      90.1090e-12
C56 34   35     25.5344e-15
L57 35   36     15.5000e-03
C58 34   36      5.0000e-12
C59 36   37    131.3387e-12
.ends
.end

