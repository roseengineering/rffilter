.SUBCKT F0 1 49
* COMMAND  : rffilter.py --g chebyshev_0.1 --bw 2500 --n 12 --l .0155 --crystal-mesh --ch 5e-12 --qu 120000 --f 8000017.0,7999933.0,7999940.0,7999945.0,7999985.0,7999996.0,8000000.0,7999991.0,7999966.0,7999945.0,7999939.0,8000026.0
* TYPE     : chebyshev_0.1
* FILTER   : crystal mesh
* ORDER    : 12
* FREQ     : 8.001743 MHz
* RE1      : 240.9
* RE2      : 240.7
* CH       : 5.0000e-12
* BW       : 2.5000e+03
* QL       : 3200.7
* QU       : 120000.0
* qo       : 37.5

* ij        q,k           TD1           TDN           CBW           Q,K      QU/QE>10
* 1      1.2055  306.9781e-06             -    2.0738e+03    3.8584e+03   31.1006e+00
* 12     0.7550  370.6146e-06    2.2652e-03    1.8874e+03  235.8743e-06   28.3049e+00
* 23     0.5644  856.1517e-06    3.0704e-03    1.4111e+03  176.3516e-06   21.1622e+00
* 34     0.5321  787.7278e-06    2.0388e-03    1.3301e+03  166.2316e-06   19.9478e+00
* 45     0.5213    1.4281e-03    2.5681e-03    1.3033e+03  162.8824e-06   19.5459e+00
* 56     0.5172    1.2116e-03    1.6336e-03    1.2929e+03  161.5758e-06   19.3891e+00
* 67     0.5160    2.0027e-03    2.0027e-03    1.2900e+03  161.2173e-06   19.3461e+00
* 78     0.5172    1.6336e-03    1.2116e-03    1.2929e+03  161.5769e-06   19.3892e+00
* 89     0.5214    2.5680e-03    1.4282e-03    1.3034e+03  162.8889e-06   19.5467e+00
* 910    0.5321    2.0388e-03  787.6913e-06    1.3302e+03  166.2327e-06   19.9479e+00
* 1011   0.5644    3.0703e-03  856.1785e-06    1.4111e+03  176.3492e-06   21.1619e+00
* 1112   0.7550    2.2653e-03  370.6053e-06    1.8874e+03  235.8779e-06   28.3054e+00
* 12     1.2055             -  306.9762e-06    2.0738e+03    3.8584e+03   31.1008e+00

* Group Delay for Lossy Q Resonators
* i         q,k           TDn            QU
* 1      1.2055  307.2958e-06  120.0000e+03
* 2      0.7550  369.7855e-06  120.0000e+03
* 3      0.5644  859.3777e-06  120.0000e+03
* 4      0.5321  783.6747e-06  120.0000e+03
* 5      0.5213    1.4405e-03  120.0000e+03
* 6      0.5172    1.2001e-03  120.0000e+03
* 7      0.5160    2.0339e-03  120.0000e+03
* -- reversed --
* i         q,k           TDn            QU
* 12     1.2055  307.2939e-06  120.0000e+03
* 11     0.7550  369.7763e-06  120.0000e+03
* 10     0.5644  859.4048e-06  120.0000e+03
* 9      0.5321  783.6383e-06  120.0000e+03
* 8      0.5214    1.4405e-03  120.0000e+03
* 7      0.5172    1.2001e-03  120.0000e+03
* 6      0.5160    2.0339e-03  120.0000e+03

* Xtal       Xtal freq     Mesh freq   Mesh offset
* 1          8000017.0     8001110.7        -632.2
* 2          7999933.0     8001738.0          -4.8
* 3          7999940.0     8001469.7        -273.1
* 4          7999945.0     8001418.7        -324.2
* 5          7999985.0     8001435.3        -307.5
* 6          7999996.0     8001437.0        -305.9
* 7          8000000.0     8001440.5        -302.3
* 8          7999991.0     8001439.9        -303.0
* 9          7999966.0     8001437.1        -305.7
* 10         7999945.0     8001473.2        -269.6
* 11         7999939.0     8001742.9          -0.0
* 12         8000026.0     8001118.3        -624.5

* Xtal              LM          LEFF     %LM Shift
* 1        15.5000e-03   18.4893e-03        19.286
* 2        15.5000e-03   18.6564e-03        20.364
* 3        15.5000e-03   18.6424e-03        20.273
* 4        15.5000e-03   18.6324e-03        20.209
* 5        15.5000e-03   18.5527e-03        19.695
* 6        15.5000e-03   18.5309e-03        19.554
* 7        15.5000e-03   18.5229e-03        19.503
* 8        15.5000e-03   18.5408e-03        19.618
* 9        15.5000e-03   18.5905e-03        19.939
* 10       15.5000e-03   18.6324e-03        20.209
* 11       15.5000e-03   18.6444e-03        20.286
* 12       15.5000e-03   18.4715e-03        19.171

* ij              CKij           CTi
* 12       90.3060e-12  135.4169e-12
* 23      120.2895e-12   17.5537e-09
* 34      127.6947e-12  310.8700e-12
* 45      130.6350e-12  262.0363e-12
* 56      132.0516e-12  277.4088e-12
* 67      132.4514e-12  279.2586e-12
* 78      132.1214e-12  282.6384e-12
* 89      130.8189e-12  281.7501e-12
* 910     127.8720e-12  278.4773e-12
* 1011    120.3621e-12  315.0820e-12
* 1112     90.3771e-12    6.3301e-03
* 1213               -  137.2074e-12

C1  1    2      25.5345e-15
L2  2    3      15.5000e-03
R3  3    4       6.4940e+00
C4  1    4       5.0000e-12
C5  4    5     135.4169e-12

C6  5    0      90.3060e-12
C7  5    6      25.5350e-15
L8  6    7      15.5000e-03
R9  7    8       6.4940e+00
C10 5    8       5.0000e-12
C11 8    9      17.5537e-09

C12 9    0     120.2895e-12
C13 9    10     25.5350e-15
L14 10   11     15.5000e-03
R15 11   12      6.4940e+00
C16 9    12      5.0000e-12
C17 12   13    310.8700e-12

C18 13   0     127.6947e-12
C19 13   14     25.5349e-15
L20 14   15     15.5000e-03
R21 15   16      6.4940e+00
C22 13   16      5.0000e-12
C23 16   17    262.0363e-12

C24 17   0     130.6350e-12
C25 17   18     25.5347e-15
L26 18   19     15.5000e-03
R27 19   20      6.4940e+00
C28 17   20      5.0000e-12
C29 20   21    277.4088e-12

C30 21   0     132.0516e-12
C31 21   22     25.5346e-15
L32 22   23     15.5000e-03
R33 23   24      6.4940e+00
C34 21   24      5.0000e-12
C35 24   25    279.2586e-12

C36 25   0     132.4514e-12
C37 25   26     25.5346e-15
L38 26   27     15.5000e-03
R39 27   28      6.4940e+00
C40 25   28      5.0000e-12
C41 28   29    282.6384e-12

C42 29   0     132.1214e-12
C43 29   30     25.5346e-15
L44 30   31     15.5000e-03
R45 31   32      6.4940e+00
C46 29   32      5.0000e-12
C47 32   33    281.7501e-12

C48 33   0     130.8189e-12
C49 33   34     25.5348e-15
L50 34   35     15.5000e-03
R51 35   36      6.4940e+00
C52 33   36      5.0000e-12
C53 36   37    278.4773e-12

C54 37   0     127.8720e-12
C55 37   38     25.5349e-15
L56 38   39     15.5000e-03
R57 39   40      6.4940e+00
C58 37   40      5.0000e-12
C59 40   41    315.0820e-12

C60 41   0     120.3621e-12
C61 41   42     25.5350e-15
L62 42   43     15.5000e-03
R63 43   44      6.4940e+00
C64 41   44      5.0000e-12
C65 44   45      6.3301e-03

C66 45   0      90.3771e-12
C67 45   46     25.5344e-15
L68 46   47     15.5000e-03
R69 47   48      6.4940e+00
C70 45   48      5.0000e-12
C71 48   49    137.2074e-12
.ends
.end

