.SUBCKT F1 1 4 5 8 9 12 13 16 17 20 21 24 25 28 29 32
* COMMAND  : rffilter.py -k chebyshev_0.5 -bw 2500 -n 8 -l 70e-3 -crystal -cp 3.7e-12 -f 5000.680e3,5000.123e3,4999.670e3,5000.235e3,5000.320e3,4999.895e3,5000.010e3,5000.485e3
* TYPE     : CHEBYSHEV_0.5
* FILTER   : CRYSTAL_MESH
* ORDER    : 8
* FREQ     : 5.001933 MHz
* RS       : 810.3
* RL       : 848.6
* BW       : 2.5000e+03
* QL       : 2000.8

* ij    qi,kij           TD0           TDn           CBW
* 01    1.7850  454.5465e-06             -    1.4006e+03
* 12    0.6580  329.4960e-06    1.2890e-03    1.6450e+03
* 23    0.5330    1.1473e-03    2.4582e-03    1.3325e+03
* 34    0.5150  682.4272e-06    1.0554e-03    1.2875e+03
* 45    0.5110    1.8509e-03    1.8172e-03    1.2775e+03
* 56    0.5150    1.0299e-03  699.3288e-06    1.2875e+03
* 67    0.5330    2.5078e-03    1.1306e-03    1.3325e+03
* 78    0.6500    1.2635e-03  337.6566e-06    1.6250e+03
* 89    1.7850             -  454.5465e-06    1.4006e+03

C1  1    2      14.4705e-15
L2  2    3      70.0000e-03
C3  1    3       3.7000e-12
C4  3    4     129.2824e-12

C5  4    0      31.2510e-12
C6  5    6      14.4737e-15
L7  6    7      70.0000e-03
C8  5    7       3.7000e-12
C9  7    8     461.1271e-09

C10 8    0      34.0121e-12
C11 9    10     14.4764e-15
L12 10   11     70.0000e-03
C13 9    11      3.7000e-12
C14 11   12     41.7101e-12

C15 12   0      35.6953e-12
C16 13   14     14.4731e-15
L17 14   15     70.0000e-03
C18 13   15      3.7000e-12
C19 15   16    312.0102e-12

C20 16   0      39.0842e-12
C21 17   18     14.4726e-15
L22 18   19     70.0000e-03
C23 17   19      3.7000e-12
C24 19   20      1.1144e-09

C25 20   0      37.1498e-12
C26 21   22     14.4751e-15
L27 22   23     70.0000e-03
C28 21   23      3.7000e-12
C29 23   24     65.3799e-12

C30 24   0      34.5333e-12
C31 25   26     14.4744e-15
L32 26   27     70.0000e-03
C33 25   27      3.7000e-12
C34 27   28    227.2237e-12

C35 28   0      30.4743e-12
C36 29   30     14.4716e-15
L37 30   31     70.0000e-03
C38 29   31      3.7000e-12
C39 31   32     70.5414e-12
.ends
.end

