.SUBCKT F1 1 10
* COMMAND: rffilter.py -g butterworth -nodal -f 10e6 -bw 400e3 -n 5 -qu 200
* TYPE:    BUTTERWORTH
* FILTER:  NODAL
* ORDER:   5
* FREQ:    10.000000 MHz 
* RS:      50.0
* RL:      50.0
* BW:      400.0000e+03
* QL:      25.0
* QU:      200.0

* ij    qi,kij           TD0           TDn           CBW
* 01    0.6180  983.6253e-09             -  647.2178e+03
* 12    1.0000    2.5752e-06    5.1503e-06  400.0018e+03
* 23    0.5559    4.1667e-06    5.1503e-06  222.3575e+03
* 34    0.5559    5.1503e-06    4.1667e-06  222.3575e+03
* 45    1.0000    5.1503e-06    2.5752e-06  400.0018e+03
* 56    0.6180             -  983.6253e-09  647.2178e+03

R1  1  2    16.1804e-03
L2  2  0    51.5040e-09
C3  1  0     4.7214e-09
C4  2  3   196.7259e-12

R5  3  4    16.1804e-03
L6  4  0    51.5040e-09
C7  3  0     4.6120e-09
C8  4  5   109.3582e-12

R9  5  6    16.1804e-03
L10 6  0    51.5040e-09
C11 5  0     4.6994e-09
C12 6  7   109.3582e-12

R13 7  8    16.1804e-03
L14 8  0    51.5040e-09
C15 7  0     4.6120e-09
C16 8  9   196.7259e-12

R17 9  10   16.1804e-03
L18 10 0    51.5040e-09
C19 9  0     4.7214e-09
.ends
.end

