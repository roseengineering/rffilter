.SUBCKT F1 1 2 3 4 5
* COMMAND  : rffilter.py -k chebyshev_0.1 -nodal -expose -f 10e6 -bw 400e3 -n 5 -qu 2000
* TYPE     : CHEBYSHEV_0.1
* FILTER   : NODAL
* ORDER    : 5
* FREQ     : 10.000000 MHz
* RS       : 50.0
* RL       : 50.0
* BW       : 400.0000e+03
* QL       : 25.0
* QU       : 2000.0

* ij    qi,kij           TD0           TDn           CBW
* 01    1.3010    2.0706e-06             -  307.4558e+03
* 12    0.7030    2.4753e-06    7.7031e-06  281.2000e+03
* 23    0.5360    5.6325e-06    4.9506e-06  214.4000e+03
* 34    0.5360    4.9506e-06    5.6325e-06  214.4000e+03
* 45    0.7030    7.7031e-06    2.4753e-06  281.2000e+03
* 56    1.3010             -    2.0706e-06  307.4558e+03

L1  1    1001   24.4666e-09
R1  1001 0     768.6395e-06
C2  1    0      10.0619e-09
C3  1    2     291.1272e-12

L4  2    1004   24.4666e-09
R4  1004 0     768.6395e-06
C5  2    0       9.8399e-09
C6  2    3     221.9689e-12

L7  3    1007   24.4666e-09
R7  1007 0     768.6395e-06
C8  3    0       9.9091e-09
C9  3    4     221.9689e-12

L10 4    1010   24.4666e-09
R10 1010 0     768.6395e-06
C11 4    0       9.8399e-09
C12 4    5     291.1272e-12

L13 5    1013   24.4666e-09
R13 1013 0     768.6395e-06
C14 5    0      10.0619e-09
.ends
.end

