.SUBCKT F0 1 2 3 4 5
* COMMAND  : rffilter.py --k chebyshev_0.1 --nodal --expose --f 10e6 --bw 400e3 --n 5 --re 50 --qu 2000
* TYPE     : chebyshev_0.1
* FILTER   : nodal
* ORDER    : 5
* FREQ     : 10.000000 MHz
* RE1      : 50.0
* RE2      : 50.0
* BW       : 400.0000e+03
* QL       : 25.0
* QU       : 2000.0
* qo       : 80.0

* ij        q,k           TD1           TDN           CBW           Q,K
* 1      1.3010    2.0706e-06             -  307.4558e+03   32.5250e+00
* 12     0.7030    2.4753e-06    7.7031e-06  281.2000e+03   28.1200e-03
* 23     0.5360    5.6325e-06    4.9506e-06  214.4000e+03   21.4400e-03
* 34     0.5360    4.9506e-06    5.6325e-06  214.4000e+03   21.4400e-03
* 45     0.7030    7.7031e-06    2.4753e-06  281.2000e+03   28.1200e-03
* 5      1.3010             -    2.0706e-06  307.4558e+03   32.5250e+00

R1  1    1001  756.1395e-06
L1  1001 0      24.0687e-09
C2  1    0      10.2282e-09
C3  1    2     295.9399e-12

R4  2    1002  756.1395e-06
L4  1002 0      24.0687e-09
C5  2    0      10.0026e-09
C6  2    3     225.6384e-12

R7  3    1003  756.1395e-06
L7  1003 0      24.0687e-09
C8  3    0      10.0729e-09
C9  3    4     225.6384e-12

R10 4    1004  756.1395e-06
L10 1004 0      24.0687e-09
C11 4    0      10.0026e-09
C12 4    5     295.9399e-12

R13 5    1005  756.1395e-06
L13 1005 0      24.0687e-09
C14 5    0      10.2282e-09
.ends
.end

